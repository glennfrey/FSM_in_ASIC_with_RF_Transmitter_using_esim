* C:\Users\glenn\eSim-Workspace\ASK\ASK.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 3/12/2022 5:03:05 PM

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U2  TX plot_v1		
v2  TX Net-_M1-Pad3_ sine		
M1  Net-_M1-Pad1_ Data Net-_M1-Pad3_ Net-_M1-Pad4_ mosfet_n		
v3  Net-_M2-Pad4_ GND DC		
M2  Net-_M1-Pad1_ Data TX Net-_M2-Pad4_ mosfet_p		
v4  GND Net-_M1-Pad4_ DC		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ ? ? Net-_U1-Pad13_ glenn_uart		
U5  Net-_U1-Pad13_ Data dac_bridge_1		
U4  GND GND GND GND GND GND GND GND Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ adc_bridge_8		
v5  Net-_U3-Pad2_ GND DC		
v1  clk GND pulse		
U6  Data plot_v1		
U3  clk Net-_U3-Pad2_ Net-_U1-Pad1_ Net-_U1-Pad2_ adc_bridge_2		
U7  clk plot_v1		

.end
