* C:\Users\glenn\eSim-Workspace\glenn_updownCounter\glenn_updownCounter.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 3/10/2022 11:01:46 PM

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U1  clk Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U1-Pad11_ glenn_updowncounter		
X1  ? ? Net-_X1-Pad3_ ? ? Net-_X1-Pad6_ Net-_U1-Pad2_ ? lm_741		
X3  Net-_U1-Pad11_ Net-_U1-Pad10_ Net-_U1-Pad9_ Net-_U1-Pad8_ Net-_U1-Pad7_ Net-_U1-Pad6_ Net-_U1-Pad5_ Net-_U1-Pad4_ GND GND Net-_X1-Pad3_ 10bitDAC		
X2  Net-_X1-Pad6_ Net-_U1-Pad2_ clk Net-_U1-Pad3_ 3_and		

.end
